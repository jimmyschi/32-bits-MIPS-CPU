----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/23/2022 09:20:47 AM
-- Design Name: 
-- Module Name: Memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Memory is
  Port (clk, reset : in std_logic;
        addr, write_data : in std_logic_vector(31 downto 0);
        MemRead, MemWrite : in std_logic;
        Mem_data : out std_logic_vector(31 downto 0)
   );
end Memory;

architecture Behavioral of Memory is
begin
process(clk,reset)
begin
    if(reset = '1') then
        Mem_data <= (others => '0');
    elsif(rising_edge(clk)) then       
      if(MemRead = '1') then
        Mem_data <= addr;
      elsif(MemWrite = '1') then
        Mem_data <= write_data;
     end if;
end if;
end process;
end Behavioral;
